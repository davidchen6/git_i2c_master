`ifndef REG_MODEL_PKG__SV
`define REG_MODEL_PKG__SV

package reg_model_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

//  `include "tb_defines.sv"

  //include sv file
//  `include "i2c_cov.sv"
  `include "reg_model.sv"

endpackage: reg_model_pkg
`endif
